`default_nettype none

module tt_um_htfab_cells (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

cell_mux cm_inst (
    .tristate_gate(uio_in[3] && ena),
    .page(ui_in[4:0]),
    .in({uio_in[2:0], ui_in[7:5]}),
    .out(uo_out)
);

assign uio_out = 0;
assign uio_oe = 0;
wire _unused = &{clk, rst_n, uio_in[7:4], 1'b0};

endmodule
